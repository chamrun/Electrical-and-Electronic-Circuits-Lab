** Profile: "SCHEMATIC1-1"  [ C:\THINGS\UNI\3RDTERM\ELEC\LAB\ELECTRICALANDELECTRONICCIRCUITSLAB\ELECLAB7\Orcad\lab7-SCHEMATIC1-1.sim ] 

** Creating circuit file "lab7-SCHEMATIC1-1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 0.1 1000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab7-SCHEMATIC1.net" 


.END
