** Profile: "SCHEMATIC1-16"  [ C:\THINGS\UNI\3RDTERM\ELEC\LAB\ELECTRICALANDELECTRONICCIRCUITSLAB\ELECLAB8\Orcad\eleclab8-SCHEMATIC1-16.sim ] 

** Creating circuit file "eleclab8-SCHEMATIC1-16.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2m 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\eleclab8-SCHEMATIC1.net" 


.END
