** Profile: "SCHEMATIC1-2"  [ C:\THINGS\UNI\3RDTERM\ELEC\LAB\ELECTRICALANDELECTRONICCIRCUITSLAB\ELECLAB8\Orcad\eleclab8-schematic1-2.sim ] 

** Creating circuit file "eleclab8-schematic1-2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 4m 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\eleclab8-SCHEMATIC1.net" 


.END
