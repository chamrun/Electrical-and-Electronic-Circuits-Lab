** Profile: "SCHEMATIC1-2"  [ C:\Things\uni\3rdTerm\Elec\Lab\ElectricalAndElectronicCircuitsLab\ElecLab7\Orcad\lab7-schematic1-2.sim ] 

** Creating circuit file "lab7-schematic1-2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20m 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab7-SCHEMATIC1.net" 


.END
