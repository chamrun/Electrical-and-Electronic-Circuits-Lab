** Profile: "SCHEMATIC1-4-2"  [ C:\THINGS\UNI\3RDTERM\ELEC\LAB\ELECTRICALANDELECTRONICCIRCUITSLAB\ELECLAB9\OrCad\lab10-schematic1-4-2.sim ] 

** Creating circuit file "lab10-schematic1-4-2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 40m 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab10-SCHEMATIC1.net" 


.END
