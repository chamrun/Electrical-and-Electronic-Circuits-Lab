** Profile: "SCHEMATIC1-3"  [ C:\Things\uni\3rdTerm\Elec\Lab\ElectricalAndElectronicCircuitsLab\ElecLab7\Orcad\lab7-SCHEMATIC1-3.sim ] 

** Creating circuit file "lab7-SCHEMATIC1-3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 1 1000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab7-SCHEMATIC1.net" 


.END
