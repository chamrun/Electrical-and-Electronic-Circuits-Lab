** Profile: "SCHEMATIC1-2-1"  [ C:\THINGS\UNI\3RDTERM\ELEC\LAB\ELECTRICALANDELECTRONICCIRCUITSLAB\ELECLAB9\OrCad\lab8-schematic1-2-1.sim ] 

** Creating circuit file "lab8-schematic1-2-1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V5 0 7 0.1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab8-SCHEMATIC1.net" 


.END
